module d_latch_mux(d,clock,q);
input d,clock;
inout q;
mux mux1(.a(q),.b(d),.s(clock),.y(q));
endmodule
