module OR_Gate(
  input A,
  input B,
  output Y);
  
  assign Y = A || B; 
  
endmodule
