module NOT_Gate(
  input A,
  output Y);
  
  assign Y = ~A; 
  
endmodule
