module inv;
  input a;
  output y;
  assign y=~a;
endmodule
